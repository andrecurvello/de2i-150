library verilog;
use verilog.vl_types.all;
entity aes_128_top_tb is
end aes_128_top_tb;
